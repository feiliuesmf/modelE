// See the end of this file for information about netcdf documentation
// and some uses in the modelE context.
//
// This template defines a netcdf file to which you can output any
// modelE variable at your choice of time frequency.
// In your customized copy of the template, you declare the
// names and dimensions of such variables.  Making these
// declarations exterior to the model streamlines the fortran
// programming but requires that you verify the consistency
// of your template with the particular model version you are using!
//
// Explanatory comments can be deleted from operational templates.
//
// Before running the model, remember to include INST_netcdf.f in
// your rundeck.
// Also, please check that your template contains no syntax errors,
// by running the 'ncgen' command:
//     ncgen your_netcdf_template
// In the absence of any errors there is no output from this command.
//
// See INST_netcdf.f concerning the fortran procedures to output your
// variables from within modelE.
//
// Netcdf output is written to the file nctemp.nc in the run directory.
// For now, this filename cannot be changed.

netcdf nctemp {

// ---------------------------------------------------------------------
dimensions:
// ---------------------------------------------------------------------
// These are example dimensions and can have any names or sizes.
// Please delete or comment out unused dimensions.
// Here, time is a record dimension allowing an unlimited
// number of timesteps to be stored in the output file.
// In contrast, hour24 would be a finite time dimension (see below).

	lon = 144 ;  // number of longitudes at 2x2.5 resolution
	lat = 90 ;   // number of latitudes  at 2x2.5 resolution
	p = 20 ;     // one possible vertical dimension
	hour24 = 24 ;  // for a moving window of hourly output
        time = UNLIMITED ; // the record dimension
// NOTE: there can only be one record dimension in a file.

// ---------------------------------------------------------------------
variables:
// ---------------------------------------------------------------------
// Replace "float" with "double" if more precision is desired.
// Please delete or comment out unused example variables.
// Attributes such as long_name, units, or missing_data can be added
// if desired.
// In the CDL notation, the order of dimensions follows the C language
// convention (the last listed dimension being most rapidly varying).
// The modelE code follows the fortran ordering convention.

// Having a record dimension, these arrays grow in size as the model runs.
	float example_ij_var(time, lat, lon) ;
	float example_ijl_var(time, p, lat, lon) ;
	float example_jl_var(time, p, lat) ;
// Note: since there can be only 1 UNLIMITED dimension in a file,
// all variables possessing this dimension should be written out
// at the same time frequency!  Otherwise, the netcdf library has
// to fill in missing values for the variables that were written
// less frequently.

// This array maintains a constant size as the model runs.
	float example_hour24_var(hour24, lat, lon) ;
// After the last hour24 index is reached, the modelE code will
// write the next data into the first hour24 index and so on.

// Special treatment to fill an entire array at once.
	float orography(lat, lon) ;
		orography:write_all = "yes" ;
// There is no requirement that variables have a time dimension.
// By default, the modelE code writes only one element of the
// most slowly varying dimension of an array as it is defined in the
// netcdf file.  To fill the entire array, an attribute write_all
// should be set to "yes" for that array, as shown here.  This behavior
// might be desired when writing out time-independent quantities such
// as orography or coordinate variables only once during a model run.

// A coordinate variable is a 1-d variable whose name is the same as
// its sole dimension.  It contains the values of that coordinate.
// Many software tools reading netcdf expect this kind of information
// to be present.
	float lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	float lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	float p(p) ;
		p:long_name = "pressure" ;
		p:units = "mb" ;

// ---------------------------------------------------------------------
data:
// ---------------------------------------------------------------------
// Here, specify the values of any coordinate variables not written to
// the output file during model initialization.  If these variables are
// to be written from the model, their write_all attribute needs to be
// set.

// 2 x 2.5 resolution
 lon = -178.75, -176.25, -173.75, -171.25, -168.75, -166.25, -163.75,
    -161.25, -158.75, -156.25, -153.75, -151.25, -148.75, -146.25, -143.75,
    -141.25, -138.75, -136.25, -133.75, -131.25, -128.75, -126.25, -123.75,
    -121.25, -118.75, -116.25, -113.75, -111.25, -108.75, -106.25, -103.75,
    -101.25, -98.75, -96.25, -93.75, -91.25, -88.75, -86.25, -83.75, -81.25,
    -78.75, -76.25, -73.75, -71.25, -68.75, -66.25, -63.75, -61.25, -58.75,
    -56.25, -53.75, -51.25, -48.75, -46.25, -43.75, -41.25, -38.75, -36.25,
    -33.75, -31.25, -28.75, -26.25, -23.75, -21.25, -18.75, -16.25, -13.75,
    -11.25, -8.75, -6.25, -3.75, -1.25, 1.25, 3.75, 6.25, 8.75, 11.25, 13.75,
    16.25, 18.75, 21.25, 23.75, 26.25, 28.75, 31.25, 33.75, 36.25, 38.75,
    41.25, 43.75, 46.25, 48.75, 51.25, 53.75, 56.25, 58.75, 61.25, 63.75,
    66.25, 68.75, 71.25, 73.75, 76.25, 78.75, 81.25, 83.75, 86.25, 88.75,
    91.25, 93.75, 96.25, 98.75, 101.25, 103.75, 106.25, 108.75, 111.25,
    113.75, 116.25, 118.75, 121.25, 123.75, 126.25, 128.75, 131.25, 133.75,
    136.25, 138.75, 141.25, 143.75, 146.25, 148.75, 151.25, 153.75, 156.25,
    158.75, 161.25, 163.75, 166.25, 168.75, 171.25, 173.75, 176.25, 178.75 ;
 lat = -89, -87, -85, -83, -81, -79, -77, -75, -73, -71, -69, -67, -65,
    -63, -61, -59, -57, -55, -53, -51, -49, -47, -45, -43, -41, -39, -37,
    -35, -33, -31, -29, -27, -25, -23, -21, -19, -17, -15, -13, -11, -9, -7,
    -5, -3, -1, 1, 3, 5, 7, 9, 11, 13, 15, 17, 19, 21, 23, 25, 27, 29, 31,
    33, 35, 37, 39, 41, 43, 45, 47, 49, 51, 53, 55, 57, 59, 61, 63, 65, 67,
    69, 71, 73, 75, 77, 79, 81, 83, 85, 87, 89 ;

}  // end of definitions

//
// See www.unidata.ucar.edu/software/netcdf for information about netcdf.
//
// More comments to be added about debugging, visualization,
// custom diagnostics, etc.
